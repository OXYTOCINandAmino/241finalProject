// stage1
module stage1
	(
		
	);
)
